`timescale 1ns/1ps
module mem_interface_tb;
// ******************************************************************
// PARAMETERS
// ******************************************************************
    parameter integer AXI_DATA_WIDTH    = 64;
    parameter integer RD_BUF_ADDR_WIDTH = 8;
    parameter integer NUM_AXI           = 4;
    parameter integer DATA_WIDTH        = 16;
    parameter integer NUM_DATA          = AXI_DATA_WIDTH*NUM_AXI/DATA_WIDTH;
    parameter integer NUM_PE            = 64;
    parameter integer VERBOSITY         = 2;
    parameter integer NAMESPACE_WIDTH   = 2;
    parameter integer TX_SIZE_WIDTH     = 10;
// ******************************************************************

// ******************************************************************
// Localparams
// ******************************************************************
    localparam integer STATE_IDLE           = 0;

    localparam integer WEIGHT_READ          = 1;
    localparam integer WEIGHT_READ_WAIT     = 2;

    localparam integer DATA_READ            = 3;
    localparam integer DATA_READ_WAIT       = 4;

    localparam integer STATE_COMPUTE        = 5;

    localparam integer WEIGHT_WRITE         = 6;
    localparam integer WEIGHT_WRITE_WAIT    = 7;

    localparam integer WEIGHT_COUNTER_WIDTH = 16;

    localparam integer WSTRB_WIDTH          = {(RD_BUF_DATA_WIDTH/8){1'b1}} * NUM_AXI;

    localparam integer RD_BUF_DATA_WIDTH    = DATA_WIDTH * NUM_DATA / NUM_AXI;
    localparam integer RD_IF_DATA_WIDTH     = DATA_WIDTH * NUM_DATA;
    localparam integer CTRL_PE_WIDTH        = (`C_LOG_2(NUM_PE/NUM_DATA) + 1) 
                                              * NUM_DATA + NAMESPACE_WIDTH;
    localparam integer SHIFTER_CTRL_WIDTH   = `C_LOG_2(NUM_DATA);
    localparam integer NUM_OPS              = 4;
    localparam integer OP_CODE_WIDTH        = `C_LOG_2 (NUM_OPS);
    localparam integer CTRL_BUF_DATA_WIDTH  = CTRL_PE_WIDTH + 
                                              SHIFTER_CTRL_WIDTH +
                                              OP_CODE_WIDTH;

    localparam integer OP_READ              = 0;
    localparam integer OP_SHIFT             = 1;
    localparam integer OP_WFI               = 2;
    localparam integer OP_WRITE             = 3;
// ******************************************************************

// ******************************************************************
// Wires and Regs
// ******************************************************************
    reg                             ACLK;
    reg                             ARESETN;
    reg                             EOI, EOC;
    wire                            compute_start;
    reg  [NUM_AXI-1:0]              axim_rvalid;
    wire [NUM_AXI-1:0]              axim_rready;
    reg  [RD_IF_DATA_WIDTH   -1:0]  axim_rdata;
    wire [RD_IF_DATA_WIDTH   -1:0]  rdata;
    wire [RD_IF_DATA_WIDTH   -1:0]  wdata;
    reg                             DATA_INOUT_WB;
    wire [CTRL_BUF_DATA_WIDTH-1:0]  ctrl_fifo_data_out;
    wire [CTRL_PE_WIDTH-1:0]        ctrl_pe;
    wire [OP_CODE_WIDTH-1:0]        ctrl_op_code;
    wire [SHIFTER_CTRL_WIDTH-1:0]   ctrl_shifter;

    wire  [RD_IF_DATA_WIDTH   -1:0]  shifter_input;
    assign shifter_input = mem_interface_tb.u_mem_if.rd_buf_data_out;

    reg                             fail_flag;

    integer                         i;
    integer                         n;

    integer                         pe_read_count_expected [ 0 : NUM_PE-1 ];
    integer                         pe_read_count_real     [ 0 : NUM_PE-1 ];
    //integer                         pe_write_count [ 0 : NUM_PE-1 ];

    wire [32*NUM_AXI-1:0]           S_AXI_ARADDR;
    wire [2*NUM_AXI-1:0]            S_AXI_ARBURST;
    wire [4*NUM_AXI-1:0]            S_AXI_ARCACHE;
    wire [6*NUM_AXI-1:0]            S_AXI_ARID;
    wire [4*NUM_AXI-1:0]            S_AXI_ARLEN;
    wire [2*NUM_AXI-1:0]            S_AXI_ARLOCK;
    wire [3*NUM_AXI-1:0]            S_AXI_ARPROT;
    wire [4*NUM_AXI-1:0]            S_AXI_ARQOS;
    wire [1*NUM_AXI-1:0]            S_AXI_ARUSER;
    wire [NUM_AXI-1:0]              S_AXI_ARREADY;
    wire [3*NUM_AXI-1:0]            S_AXI_ARSIZE;
    wire [NUM_AXI-1:0]              S_AXI_ARVALID;
    wire [32*NUM_AXI-1:0]           S_AXI_AWADDR;
    wire [2*NUM_AXI-1:0]            S_AXI_AWBURST;
    wire [4*NUM_AXI-1:0]            S_AXI_AWCACHE;
    wire [6*NUM_AXI-1:0]            S_AXI_AWID;
    wire [4*NUM_AXI-1:0]            S_AXI_AWLEN;
    wire [2*NUM_AXI-1:0]            S_AXI_AWLOCK;
    wire [3*NUM_AXI-1:0]            S_AXI_AWPROT;
    wire [4*NUM_AXI-1:0]            S_AXI_AWQOS;
    wire [1*NUM_AXI-1:0]            S_AXI_AWUSER;
    wire [NUM_AXI-1:0]              S_AXI_AWREADY;
    wire [3*NUM_AXI-1:0]            S_AXI_AWSIZE;
    wire [NUM_AXI-1:0]              S_AXI_AWVALID;
    wire [6*NUM_AXI-1:0]            S_AXI_BID;
    wire [1*NUM_AXI-1:0]            S_AXI_BUSER;
    wire [NUM_AXI-1:0]              S_AXI_BREADY;
    wire [2*NUM_AXI-1:0]            S_AXI_BRESP;
    wire [NUM_AXI-1:0]              S_AXI_BVALID;
    wire [RD_IF_DATA_WIDTH-1:0]     S_AXI_RDATA;
    wire [6*NUM_AXI-1:0]            S_AXI_RID;
    wire [1*NUM_AXI-1:0]            S_AXI_RUSER;
    wire [NUM_AXI-1:0]              S_AXI_RLAST;
    wire [NUM_AXI-1:0]              S_AXI_RREADY;
    wire [2*NUM_AXI-1:0]            S_AXI_RRESP;
    wire [NUM_AXI-1:0]              S_AXI_RVALID;
    wire [RD_IF_DATA_WIDTH-1:0]     S_AXI_WDATA;
    wire [6*NUM_AXI-1:0]            S_AXI_WID;
    wire [1*NUM_AXI-1:0]            S_AXI_WUSER;
    wire [NUM_AXI-1:0]              S_AXI_WLAST;
    wire [NUM_AXI-1:0]              S_AXI_WREADY;
    wire [WSTRB_WIDTH-1:0]          S_AXI_WSTRB;
    wire [NUM_AXI-1:0]              S_AXI_WVALID;

    // WRITE from BRAM to DDR
    wire [NUM_AXI-1:0]              outBuf_empty;
    wire [NUM_AXI-1:0]              outBuf_pop;
    wire [RD_IF_DATA_WIDTH-1:0]     data_from_outBuf;

    // READ from DDR to BRAM
    wire [RD_IF_DATA_WIDTH-1:0]     data_to_inBuf;
    wire [NUM_AXI-1:0]              inBuf_push;
    wire [NUM_AXI-1:0]              inBuf_full;

    // TXN REQ
    wire [NUM_AXI-1:0]              rx_req;
    wire [NUM_AXI*TX_SIZE_WIDTH-1:0]rx_req_size;
    wire [NUM_AXI-1:0]              rx_done;
    wire [NUM_AXI*32-1:0]           rx_addr;

    reg                             start;

    reg  [RD_IF_DATA_WIDTH-1:0]   expected_data_ram [0:4095];
// ******************************************************************

// ******************************************************************
// AXI Master driver
// ******************************************************************
genvar gen;
for (gen=0; gen<NUM_AXI; gen=gen+1)
begin : AXI_DRIVERS
    localparam integer wstrb_width = RD_BUF_DATA_WIDTH/8;
    axi_master_tb_driver
    #(
        .C_M_AXI_DATA_WIDTH         ( RD_BUF_DATA_WIDTH         ),
        .DATA_WIDTH                 ( DATA_WIDTH                ),
        .TX_SIZE_WIDTH              ( TX_SIZE_WIDTH             )
    ) u_axim_driver (
        .ACLK                       ( ACLK                      ),
        .ARESETN                    ( ARESETN                   ),
        .M_AXI_AWID                 ( S_AXI_AWID[6*gen+:6]      ),
        .M_AXI_AWADDR               ( S_AXI_AWADDR[32*gen+:32]  ),
        .M_AXI_AWLEN                ( S_AXI_AWLEN[4*gen+:4]     ),
        .M_AXI_AWSIZE               ( S_AXI_AWSIZE[3*gen+:3]    ),
        .M_AXI_AWBURST              ( S_AXI_AWBURST[2*gen+:2]   ),
        .M_AXI_AWLOCK               ( S_AXI_AWLOCK[2*gen+:2]    ),
        .M_AXI_AWCACHE              ( S_AXI_AWCACHE[4*gen+:4]   ),
        .M_AXI_AWPROT               ( S_AXI_AWPROT[3*gen+:3]    ),
        .M_AXI_AWQOS                ( S_AXI_AWQOS[4*gen+:4]     ),
        .M_AXI_AWUSER               ( S_AXI_AWUSER[gen+:1]      ),
        .M_AXI_AWVALID              ( S_AXI_AWVALID[gen+:1]     ),
        .M_AXI_AWREADY              ( S_AXI_AWREADY[gen+:1]     ),
        .M_AXI_WID                  ( S_AXI_WID[6*gen+:6]       ),
        .M_AXI_WDATA                ( S_AXI_WDATA[RD_BUF_DATA_WIDTH*gen+:RD_BUF_DATA_WIDTH]               ),
        .M_AXI_WSTRB                ( S_AXI_WSTRB[wstrb_width*gen+:wstrb_width]               ),
        .M_AXI_WLAST                ( S_AXI_WLAST[gen+:1]       ),
        .M_AXI_WUSER                ( S_AXI_WUSER[gen+:1]       ),
        .M_AXI_WVALID               ( S_AXI_WVALID[gen+:1]      ),
        .M_AXI_WREADY               ( S_AXI_WREADY[gen+:1]      ),
        .M_AXI_BID                  ( S_AXI_BID[6*gen+:6]       ),
        .M_AXI_BRESP                ( S_AXI_BRESP[2*gen+:2]     ),
        .M_AXI_BUSER                ( S_AXI_BUSER[gen+:1]       ),
        .M_AXI_BVALID               ( S_AXI_BVALID[gen+:1]      ),
        .M_AXI_BREADY               ( S_AXI_BREADY[gen+:1]      ),
        .M_AXI_ARID                 ( S_AXI_ARID[6*gen+:6]      ),
        .M_AXI_ARADDR               ( S_AXI_ARADDR[32*gen+:32]  ),
        .M_AXI_ARLEN                ( S_AXI_ARLEN[4*gen+:4]     ),
        .M_AXI_ARSIZE               ( S_AXI_ARSIZE[3*gen+:3]    ),
        .M_AXI_ARBURST              ( S_AXI_ARBURST[2*gen+:2]   ),
        .M_AXI_ARLOCK               ( S_AXI_ARLOCK[2*gen+:2]    ),
        .M_AXI_ARCACHE              ( S_AXI_ARCACHE[4*gen+:4]   ),
        .M_AXI_ARPROT               ( S_AXI_ARPROT[3*gen+:3]    ),
        .M_AXI_ARQOS                ( S_AXI_ARQOS[4*gen+:4]     ),
        .M_AXI_ARUSER               ( S_AXI_ARUSER[gen+:1]      ),
        .M_AXI_ARVALID              ( S_AXI_ARVALID[gen+:1]     ),
        .M_AXI_ARREADY              ( S_AXI_ARREADY[gen+:1]     ),
        .M_AXI_RID                  ( S_AXI_RID[6*gen+:6]       ),
        .M_AXI_RDATA                ( S_AXI_RDATA[RD_BUF_DATA_WIDTH*gen+:RD_BUF_DATA_WIDTH]               ),
        .M_AXI_RRESP                ( S_AXI_RRESP[2*gen+:2]     ),
        .M_AXI_RLAST                ( S_AXI_RLAST[gen+:1]       ),
        .M_AXI_RUSER                ( S_AXI_RUSER[gen+:1]       ),
        .M_AXI_RVALID               ( S_AXI_RVALID[gen+:1]      ),
        .M_AXI_RREADY               ( S_AXI_RREADY[gen+:1]      ),
        .outBuf_empty               ( outBuf_empty[gen+:1]      ),
        .outBuf_pop                 ( outBuf_pop[gen+:1]        ),
        .data_from_outBuf           ( data_from_outBuf[RD_BUF_DATA_WIDTH*gen+:RD_BUF_DATA_WIDTH]          ),
        .data_to_inBuf              ( data_to_inBuf[RD_BUF_DATA_WIDTH*gen+:RD_BUF_DATA_WIDTH]             ),
        .inBuf_push                 ( inBuf_push[gen+:1]        ),
        .inBuf_full                 ( inBuf_full[gen+:1]        ),
        .rx_req                     ( rx_req[gen+:1]            ),
        .rx_req_size                ( rx_req_size[TX_SIZE_WIDTH*gen+:TX_SIZE_WIDTH]               ),
        .rx_addr                    ( rx_addr[gen*32+:32]                   ),
        .rx_done                    ( rx_done[gen]           )
    );
end
// ******************************************************************

// ******************************************************************
// DUT - MEM Interface
// ******************************************************************
  mem_interface #(
    .DATA_WIDTH             ( DATA_WIDTH            ),
    .RD_BUF_ADDR_WIDTH      ( RD_BUF_ADDR_WIDTH     ),
    .NUM_DATA               ( NUM_DATA              ),
    .NUM_PE                 ( NUM_PE                ),
    .NUM_AXI                ( NUM_AXI               ),
    .TX_SIZE_WIDTH          ( TX_SIZE_WIDTH         )
  ) u_mem_if (
    .ACLK                   ( ACLK                  ), //input
    .ARESETN                ( ARESETN               ), //input
    .compute_start          ( compute_start         ), //output
    .rdata                  ( rdata                 ), //input
    .wdata                  ( wdata                 ), //output
    .DATA_INOUT_WB          ( DATA_INOUT_WB         ), //input
    .EOI                    ( EOI                   ), //input
    .EOC                    ( EOC                   ), //input
    .CTRL_PE                ( ctrl_pe               ), //output
    .start                  ( start                 ), //input
    .DATA_IO_DIR            ( DATA_IO_DIR           ), //output

    .S_AXI_ARADDR           ( S_AXI_ARADDR          ), //output
    .S_AXI_ARBURST          ( S_AXI_ARBURST         ), //output
    .S_AXI_ARCACHE          ( S_AXI_ARCACHE         ), //output
    .S_AXI_ARID             ( S_AXI_ARID            ), //output
    .S_AXI_ARLEN            ( S_AXI_ARLEN           ), //output
    .S_AXI_ARLOCK           ( S_AXI_ARLOCK          ), //output
    .S_AXI_ARPROT           ( S_AXI_ARPROT          ), //output
    .S_AXI_ARQOS            ( S_AXI_ARQOS           ), //output
    .S_AXI_ARUSER           ( S_AXI_ARUSER          ), //output
    .S_AXI_ARREADY          ( S_AXI_ARREADY         ), //input
    .S_AXI_ARSIZE           ( S_AXI_ARSIZE          ), //output
    .S_AXI_ARVALID          ( S_AXI_ARVALID         ), //output
    .S_AXI_AWADDR           ( S_AXI_AWADDR          ), //output
    .S_AXI_AWBURST          ( S_AXI_AWBURST         ), //output
    .S_AXI_AWCACHE          ( S_AXI_AWCACHE         ), //output
    .S_AXI_AWID             ( S_AXI_AWID            ), //output
    .S_AXI_AWLEN            ( S_AXI_AWLEN           ), //output
    .S_AXI_AWLOCK           ( S_AXI_AWLOCK          ), //output
    .S_AXI_AWPROT           ( S_AXI_AWPROT          ), //output
    .S_AXI_AWQOS            ( S_AXI_AWQOS           ), //output
    .S_AXI_AWUSER           ( S_AXI_AWUSER          ), //output
    .S_AXI_AWREADY          ( S_AXI_AWREADY         ), //input
    .S_AXI_AWSIZE           ( S_AXI_AWSIZE          ), //output
    .S_AXI_AWVALID          ( S_AXI_AWVALID         ), //output
    .S_AXI_BID              ( S_AXI_BID             ), //input
    .S_AXI_BUSER            ( S_AXI_BUSER           ), //input
    .S_AXI_BREADY           ( S_AXI_BREADY          ), //output
    .S_AXI_BRESP            ( S_AXI_BRESP           ), //input
    .S_AXI_BVALID           ( S_AXI_BVALID          ), //input
    .S_AXI_RDATA            ( S_AXI_RDATA           ), //input
    .S_AXI_RID              ( S_AXI_RID             ), //input
    .S_AXI_RUSER            ( S_AXI_RUSER           ), //input
    .S_AXI_RLAST            ( S_AXI_RLAST           ), //input
    .S_AXI_RREADY           ( S_AXI_RREADY          ), //output
    .S_AXI_RRESP            ( S_AXI_RRESP           ), //input
    .S_AXI_RVALID           ( S_AXI_RVALID          ), //input
    .S_AXI_WDATA            ( S_AXI_WDATA           ), //output
    .S_AXI_WID              ( S_AXI_WID             ), //output
    .S_AXI_WUSER            ( S_AXI_WUSER           ), //output
    .S_AXI_WLAST            ( S_AXI_WLAST           ), //output
    .S_AXI_WREADY           ( S_AXI_WREADY          ), //input
    .S_AXI_WSTRB            ( S_AXI_WSTRB           ), //output
    .S_AXI_WVALID           ( S_AXI_WVALID          )  //output

    //.rx_req                 ( rx_req                ), //input
    //.rx_req_size            ( rx_req_size           ), //input
    //.rx_done                ( rx_done               ), //output
    //.rx_addr                ( rx_addr               )  //input
  );
// ******************************************************************


//--------------------------------------------------------------------------------------
task test_main;
    begin
        repeat(20) begin
            AXI_DRIVERS[0].u_axim_driver.request_random_tx;
            $display ("AXI 0 done");
            AXI_DRIVERS[1].u_axim_driver.request_random_tx;
            $display ("AXI 1 done");
            AXI_DRIVERS[2].u_axim_driver.request_random_tx;
            $display ("AXI 2 done");
            AXI_DRIVERS[3].u_axim_driver.request_random_tx;
            $display ("AXI 3 done");
        end
        AXI_DRIVERS[0].u_axim_driver.check_fail;
        AXI_DRIVERS[1].u_axim_driver.check_fail;
        AXI_DRIVERS[2].u_axim_driver.check_fail;
        AXI_DRIVERS[3].u_axim_driver.check_fail;
        //AXI_DRIVERS[0].u_axim_driver.test_pass;
    end
endtask
//--------------------------------------------------------------------------------------

//--------------------------------------------------------------------------------------
wire ctrl_buf_rd_en       = mem_interface_tb.u_mem_if.u_if_controller.ctrl_buf_read_en;
reg ctrl_buf_rd_en_reg;
wire [11:0] ctrl_buf_addr = mem_interface_tb.u_mem_if.u_if_controller.ctrl_buf_addr;
assign ctrl_fifo_data_out = mem_interface_tb.u_mem_if.u_if_controller.ctrl_buf_data_out;

wire [NUM_AXI*RD_BUF_ADDR_WIDTH-1:0] rd_address_received;

generate
for(gen=0; gen<NUM_AXI; gen=gen+1)
begin
    assign rd_address_received[gen*RD_BUF_ADDR_WIDTH+:RD_BUF_ADDR_WIDTH] = mem_interface_tb.u_mem_if.AXI_RD_BUF[gen].read_buffer.rd_pointer;
end
endgenerate

integer num_instructions;
initial begin
  num_instructions = 0;
end

always @(posedge ACLK)
begin
  if (ctrl_buf_rd_en)
    num_instructions = num_instructions + 1;
end

//--------------------------------------------------------------------------------------
task rand_instruction;
  input integer num_ins;
  reg  [CTRL_PE_WIDTH-1:0]        ctrl_pe;
  reg  [OP_CODE_WIDTH-1:0]        ctrl_op_code;
  reg  [SHIFTER_CTRL_WIDTH-1:0]   ctrl_shifter;
  reg  [CTRL_BUF_DATA_WIDTH-1:0]  ctrl_buf_data_in;
  reg  [DATA_WIDTH-1:0]           rd_data_addr;
  integer                         expected_data_addr;
  reg  [RD_IF_DATA_WIDTH-1:0]     tmp;
  integer n, m, pe_id;
  begin
    expected_data_addr = 0;
    rd_data_addr = 0;
    for (n=0; n<NUM_PE; n=n+1)
    begin
      pe_read_count_expected[n] = 0;
      pe_read_count_real[n] = 0;
      //pe_write_count[n] = 0;
    end
    for (n=0; n<num_ins; n=n+1)
    begin
      if (n > 0)
      begin
        ctrl_pe       = {$random, $random};
        ctrl_op_code  = {$random, $random} % 3;
        ctrl_shifter  = {$random, $random};
        case (ctrl_op_code)
          0:begin
            rd_data_addr = rd_data_addr + 1;
          end
          1:begin
            tmp = {
              (rd_data_addr << 2) + 2'h3, 
              (rd_data_addr << 2) + 2'h2, 
              (rd_data_addr << 2) + 2'h1, 
              (rd_data_addr << 2) + 2'h0,
              (rd_data_addr << 2) + 2'h3, 
              (rd_data_addr << 2) + 2'h2, 
              (rd_data_addr << 2) + 2'h1, 
              (rd_data_addr << 2) + 2'h0,
              (rd_data_addr << 2) + 2'h3, 
              (rd_data_addr << 2) + 2'h2, 
              (rd_data_addr << 2) + 2'h1, 
              (rd_data_addr << 2) + 2'h0,
              (rd_data_addr << 2) + 2'h3, 
              (rd_data_addr << 2) + 2'h2, 
              (rd_data_addr << 2) + 2'h1, 
              (rd_data_addr << 2) + 2'h0
              };
            expected_data_ram[expected_data_addr] = {tmp, tmp, tmp} >> ctrl_shifter*DATA_WIDTH;
            $display ("Expected Data : %h", expected_data_ram[expected_data_addr]);
            expected_data_addr = expected_data_addr + 1;
          end
          default:begin
          end
        endcase
      end
      else begin
        ctrl_pe       = {$random, $random};
        ctrl_op_code  = 0;
        ctrl_shifter  = {$random, $random};
      end
      if (VERBOSITY > 2) $display ("ADDR: %h, OP_CODE = %h", n, ctrl_op_code);
      for (m=0; m<NUM_DATA; m=m+1)
      begin
        if (ctrl_pe[NAMESPACE_WIDTH+(3)*m+:1] && ctrl_op_code == 1)
        begin
          pe_id = (m<<2)+ctrl_pe[NAMESPACE_WIDTH+(3)*m+1+:2];
          if (VERBOSITY > 2) $display ("Lane %d, PE_ID %d", m, pe_id);
          pe_read_count_expected[pe_id] = pe_read_count_expected[pe_id] + 1;
        end
      end
      ctrl_pe[NAMESPACE_WIDTH-1:0] = `NAMESPACE_MEM_DATA;
      ctrl_buf_data_in = {ctrl_pe, ctrl_op_code, ctrl_shifter};
      mem_interface_tb.u_mem_if.u_if_controller.u_ctrl_buf.mem[n] = ctrl_buf_data_in;
    end
    ctrl_pe       = {$random, $random};
    ctrl_op_code  = 2;
    ctrl_shifter  = {$random, $random};
    ctrl_pe[NAMESPACE_WIDTH-1:0] = `NAMESPACE_MEM_DATA;
    ctrl_buf_data_in = {ctrl_pe, ctrl_op_code, ctrl_shifter};
    mem_interface_tb.u_mem_if.u_if_controller.u_ctrl_buf.mem[num_ins] = ctrl_buf_data_in;
  end
endtask
//--------------------------------------------------------------------------------------

//--------------------------------------------------------------------------------------
task check_fail;
    if (fail_flag && ARESETN) 
    begin
        $display("%c[1;31m",27);
        $display ("Test Failed");
        $display("%c[0m",27);
        @(posedge ACLK);
        @(posedge ACLK);
        $finish;
    end
endtask
//--------------------------------------------------------------------------------------

// ******************************************************************
// TestBench
// ******************************************************************
initial
begin
    $dumpfile("hw-imp/bin/waveform/mem_interface.vcd");
    $dumpvars(0,mem_interface_tb);
end

initial 
begin
  $display("***************************************");
  $display ("Testing Read IF");
  $display("***************************************");
  n = 0;
  DATA_INOUT_WB = 1;
  ACLK = 0;
  ARESETN = 1;
  @(negedge ACLK);
  ARESETN = 0;
  set_weight_reads;
  @(negedge ACLK);
  ARESETN = 1;

  @(negedge ACLK);

  //test_main;

  //$display("%c[1;32m",27);
  //$display ("Test Passed");
  //$display("%c[0m",27);

  //#10000;
  //check_fail;
  //$finish;
end

initial begin
  EOI = 0;
  EOC = 0;
  wait (ARESETN);
  start = 1;
end

wire [2:0] state = mem_interface_tb.u_mem_if.u_if_controller.state;
reg [16-1:0] a;
integer pe_id_count;
initial
begin
  rand_instruction(100);
  $display ("Testing random instructions");
  wait(num_instructions == 100);
  wait (state == 0);
  for (pe_id_count = 0; pe_id_count < NUM_PE; pe_id_count = pe_id_count + 1)
  begin
    if (pe_read_count_expected[pe_id_count] !== pe_read_count_real[pe_id_count]) begin
      fail_flag = 1;
    end
  end
  @(negedge ACLK);
  check_fail;

  check_weight_reads;
  check_fail;

  $display("%c[1;32m",27);
  $display ("**************************************************");
  $display ("Test Passed");
  $display ("**************************************************");
  $display("%c[0m",27);
  $finish;
end

task check_weight_reads;
  begin
    for (pe_id_count = 0; pe_id_count < NUM_PE; pe_id_count = pe_id_count + 1)
    begin
      a = (mem_interface_tb.u_mem_if.u_if_controller.counter_init[pe_id_count >> 2] >> (16*(pe_id_count%4))) & 64'hFFFF;
      if (weight_read_count[pe_id_count] !== a)
      begin
        $display ("PE_ID = %d, Weight Reads = %d, Expected Weight Reads = %d", 
          pe_id_count, weight_read_count[pe_id_count], a);
        fail_flag = 1;
        check_fail;
      end
    end
  end
endtask

always #1 ACLK = ~ACLK;

always @ (posedge ACLK)
begin
  check_fail;
  DATA_INOUT_WB = $random;
end

wire shifter_rd_en = mem_interface_tb.u_mem_if.shifter_rd_en;
integer addr;
initial begin
  addr = 0;
end
always @(posedge ACLK)
begin
  if (shifter_rd_en)
    check_shifter_output;
end

task check_shifter_output;
  integer n, m, pe_id;
  reg valid;
  reg [1:0] namespace;
  begin
    // for (n=0; n<NUM_DATA; n=n+1)
    // begin
    //   pe_id = (n<<2)+ctrl_pe[NAMESPACE_WIDTH+(3)*n+1+:2];
    //   valid = ctrl_pe[NAMESPACE_WIDTH+(3)*n+:1];
    //   if (valid) $display ("state = %d PE ID = %d", state, pe_id);
    // end
    namespace = ctrl_pe[NAMESPACE_WIDTH-1:0];
    @(negedge ACLK);
    if (wdata !== expected_data_ram[addr] && namespace == `NAMESPACE_MEM_DATA) begin
      $display ("Got Data      : %h", wdata);
      $display ("Expected Data : %h", expected_data_ram[addr]);
      fail_flag = 1;
    end
    else if (VERBOSITY > 2) begin
      $display ("Got Data      : %h", wdata);
      $display ("Expected Data : %h", expected_data_ram[addr]);
    end
    if (namespace == `NAMESPACE_MEM_DATA) addr = addr + 1;
    // for (n=0; n<NUM_DATA; n=n+1)
    // begin
    //   pe_id = (n<<2)+ctrl_pe[NAMESPACE_WIDTH+(3)*n+1+:2];
    //   valid = ctrl_pe[NAMESPACE_WIDTH+(3)*n+:1];
    //   if (valid) $display ("state = %d PE ID = %d", state, pe_id);
    // end
  end
endtask

always @(posedge ACLK)
begin
  count_pe_reads;
end

task count_pe_reads;
  integer n, m, pe_id;
  reg valid;
  reg [1:0] namespace;
  if (ctrl_pe[NAMESPACE_WIDTH-1:0] == `NAMESPACE_MEM_DATA)
  begin
    if (VERBOSITY > 2) $display ("--");
    for (n=0; n<NUM_DATA; n=n+1)
    begin
      pe_id = (n<<2)+ctrl_pe[NAMESPACE_WIDTH+(3)*n+1+:2];
      valid = ctrl_pe[NAMESPACE_WIDTH+(3)*n+:1];
      if (valid) begin
        pe_read_count_real[pe_id] = pe_read_count_real[pe_id] + 1;
        if (VERBOSITY > 2) $display ("PE_ID - %d, Expected Reads = %d, Actual = %d",
          pe_id, pe_read_count_expected[pe_id], pe_read_count_real[pe_id]);
      end
    end
    if (VERBOSITY > 2) $display ("--");
  end
endtask

always @(posedge ACLK)
begin
  if (compute_start)
    compute;
end

task compute;
  begin
    repeat (10) @(negedge ACLK);
    if (num_instructions < 101) begin
      EOI = 1;
      EOC = 0;
    end
    else begin
      EOI = 0;
      EOC = 1;
    end
    @(negedge ACLK);
      EOI = 0;
      EOC = 0;
  end
endtask

integer weight_read_count [ NUM_PE-1 : 0 ];

initial begin
end

always @(posedge ACLK)
begin
  if (ARESETN == 0 || (shifter_rd_en && ctrl_pe[NAMESPACE_WIDTH-1:0] == `NAMESPACE_MEM_WEIGHT && DATA_IO_DIR == 0))
  begin
    count_weight_reads;
  end
end

task set_weight_reads;
  begin
    for (i=0; i<NUM_PE; i=i+1)
    begin
      //mem_interface_tb.u_mem_if.u_if_controller.counter_init[i] = {16'd16, 16'd9, 16'd6, 16'd8};
      mem_interface_tb.u_mem_if.u_if_controller.counter_init[i] = {$random & 32'h00FF00FF, $random & 32'h00FF00FF};
    end
  end
endtask

task count_weight_reads;
  integer n, pe_id;
  reg valid;
  begin
    if (ARESETN == 0)
    begin
      for (n=0; n<NUM_PE; n=n+1)
      begin
        weight_read_count[n] = 0;
      end
    end
    for (n=0; n<NUM_DATA; n=n+1)
    begin
      pe_id = (n<<2)+ctrl_pe[NAMESPACE_WIDTH+(3)*n+1+:2];
      valid = ctrl_pe[NAMESPACE_WIDTH+(3)*n+:1];
      if (valid)
      begin
        weight_read_count[pe_id] = weight_read_count[pe_id] + 1;
      end
    end
  end
endtask

// ******************************************************************

endmodule
