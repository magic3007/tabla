`timescale 1ns / 100ps

//INDEXES FOR EACH NAMESPACE
`define INDEX_INST 		6
`define INDEX_DATA 		6
`define INDEX_WEIGHT 	6
`define INDEX_META 		2
`define INDEX_INTERIM 2


//NUMBER OF VALID PEs
`define NUM_PE_VALID 6

//COMPUTE ELEMENTS
//`define GAUSSIAN
//`define DIV
//`define SQRT
`define SIGMOID


