`timescale 1ns/1ps
module sigmoid (
    in,
    out
);
    //--------------------------------------------------------------------------------------
    //parameter LEN  = 9;
    //parameter OUTLEN = 7;
    parameter LEN = 32;
    parameter FRACTION = 15;

    //--------------------------------------------------------------------------------------
    input[LEN - 1: 0]   in;
    output[LEN - 1: 0] out;
    reg[LEN - 1: 0] res;
    wire[6:0] index;

    assign out = res;
    always @(index)
    begin
        case(index) //128 lut entries here
            7'd0: res = 32'b00000000000000000100000010000000; // input=0.015625, output=0.503906170529
            7'd1: res = 32'b00000000000000000100000110000000; // input=0.046875, output=0.511716604704
            7'd2: res = 32'b00000000000000000100001010000000; // input=0.078125, output=0.519521321952
            7'd3: res = 32'b00000000000000000100001101111111; // input=0.109375, output=0.52731652338
            7'd4: res = 32'b00000000000000000100010001111110; // input=0.140625, output=0.535098428627
            7'd5: res = 32'b00000000000000000100010101111101; // input=0.171875, output=0.542863283173
            7'd6: res = 32'b00000000000000000100011001111010; // input=0.203125, output=0.550607365535
            7'd7: res = 32'b00000000000000000100011101110111; // input=0.234375, output=0.558326994335
            7'd8: res = 32'b00000000000000000100100001110011; // input=0.265625, output=0.566018535196
            7'd9: res = 32'b00000000000000000100100101101110; // input=0.296875, output=0.573678407453
            7'd10: res = 32'b00000000000000000100101001101000; // input=0.328125, output=0.581303090644
            7'd11: res = 32'b00000000000000000100101101100001; // input=0.359375, output=0.588889130768
            7'd12: res = 32'b00000000000000000100110001011000; // input=0.390625, output=0.596433146265
            7'd13: res = 32'b00000000000000000100110101001110; // input=0.421875, output=0.603931833726
            7'd14: res = 32'b00000000000000000100111001000010; // input=0.453125, output=0.611381973294
            7'd15: res = 32'b00000000000000000100111100110100; // input=0.484375, output=0.618780433744
            7'd16: res = 32'b00000000000000000101000000100101; // input=0.515625, output=0.626124177228
            7'd17: res = 32'b00000000000000000101000100010100; // input=0.546875, output=0.633410263678
            7'd18: res = 32'b00000000000000000101001000000000; // input=0.578125, output=0.64063585484
            7'd19: res = 32'b00000000000000000101001011101011; // input=0.609375, output=0.647798217952
            7'd20: res = 32'b00000000000000000101001111010100; // input=0.640625, output=0.654894729042
            7'd21: res = 32'b00000000000000000101010010111010; // input=0.671875, output=0.66192287585
            7'd22: res = 32'b00000000000000000101010110011110; // input=0.703125, output=0.668880260371
            7'd23: res = 32'b00000000000000000101011001111111; // input=0.734375, output=0.675764601019
            7'd24: res = 32'b00000000000000000101011101011111; // input=0.765625, output=0.682573734412
            7'd25: res = 32'b00000000000000000101100000111011; // input=0.796875, output=0.689305616785
            7'd26: res = 32'b00000000000000000101100100010101; // input=0.828125, output=0.695958325033
            7'd27: res = 32'b00000000000000000101100111101101; // input=0.859375, output=0.702530057395
            7'd28: res = 32'b00000000000000000101101011000001; // input=0.890625, output=0.709019133785
            7'd29: res = 32'b00000000000000000101101110010011; // input=0.921875, output=0.715423995783
            7'd30: res = 32'b00000000000000000101110001100010; // input=0.953125, output=0.721743206298
            7'd31: res = 32'b00000000000000000101110100101110; // input=0.984375, output=0.727975448906
            7'd32: res = 32'b00000000000000000101110111111000; // input=1.015625, output=0.7341195269
            7'd33: res = 32'b00000000000000000101111010111110; // input=1.046875, output=0.740174362039
            7'd34: res = 32'b00000000000000000101111110000001; // input=1.078125, output=0.746138993031
            7'd35: res = 32'b00000000000000000110000001000010; // input=1.109375, output=0.75201257376
            7'd36: res = 32'b00000000000000000110000011111111; // input=1.140625, output=0.757794371275
            7'd37: res = 32'b00000000000000000110000110111010; // input=1.171875, output=0.763483763554
            7'd38: res = 32'b00000000000000000110001001110001; // input=1.203125, output=0.769080237071
            7'd39: res = 32'b00000000000000000110001100100110; // input=1.234375, output=0.774583384165
            7'd40: res = 32'b00000000000000000110001111010111; // input=1.265625, output=0.779992900254
            7'd41: res = 32'b00000000000000000110010010000101; // input=1.296875, output=0.785308580888
            7'd42: res = 32'b00000000000000000110010100110000; // input=1.328125, output=0.79053031867
            7'd43: res = 32'b00000000000000000110010111011000; // input=1.359375, output=0.795658100063
            7'd44: res = 32'b00000000000000000110011001111101; // input=1.390625, output=0.800692002096
            7'd45: res = 32'b00000000000000000110011100011111; // input=1.421875, output=0.805632188981
            7'd46: res = 32'b00000000000000000110011110111110; // input=1.453125, output=0.81047890867
            7'd47: res = 32'b00000000000000000110100001011010; // input=1.484375, output=0.815232489352
            7'd48: res = 32'b00000000000000000110100011110010; // input=1.515625, output=0.819893335914
            7'd49: res = 32'b00000000000000000110100110001000; // input=1.546875, output=0.824461926377
            7'd50: res = 32'b00000000000000000110101000011011; // input=1.578125, output=0.828938808321
            7'd51: res = 32'b00000000000000000110101010101010; // input=1.609375, output=0.833324595312
            7'd52: res = 32'b00000000000000000110101100110111; // input=1.640625, output=0.837619963333
            7'd53: res = 32'b00000000000000000110101111000001; // input=1.671875, output=0.841825647252
            7'd54: res = 32'b00000000000000000110110001001000; // input=1.703125, output=0.845942437309
            7'd55: res = 32'b00000000000000000110110011001100; // input=1.734375, output=0.849971175658
            7'd56: res = 32'b00000000000000000110110101001101; // input=1.765625, output=0.853912752952
            7'd57: res = 32'b00000000000000000110110111001011; // input=1.796875, output=0.85776810499
            7'd58: res = 32'b00000000000000000110111001000111; // input=1.828125, output=0.861538209431
            7'd59: res = 32'b00000000000000000110111011000000; // input=1.859375, output=0.865224082577
            7'd60: res = 32'b00000000000000000110111100110110; // input=1.890625, output=0.868826776238
            7'd61: res = 32'b00000000000000000110111110101001; // input=1.921875, output=0.872347374678
            7'd62: res = 32'b00000000000000000111000000011010; // input=1.953125, output=0.875786991648
            7'd63: res = 32'b00000000000000000111000010001000; // input=1.984375, output=0.87914676751
            7'd64: res = 32'b00000000000000000011111110000000; // input=-0.015625, output=0.496093829471
            7'd65: res = 32'b00000000000000000011111010000000; // input=-0.046875, output=0.488283395296
            7'd66: res = 32'b00000000000000000011110110000000; // input=-0.078125, output=0.480478678048
            7'd67: res = 32'b00000000000000000011110010000001; // input=-0.109375, output=0.47268347662
            7'd68: res = 32'b00000000000000000011101110000010; // input=-0.140625, output=0.464901571373
            7'd69: res = 32'b00000000000000000011101010000011; // input=-0.171875, output=0.457136716827
            7'd70: res = 32'b00000000000000000011100110000110; // input=-0.203125, output=0.449392634465
            7'd71: res = 32'b00000000000000000011100010001001; // input=-0.234375, output=0.441673005665
            7'd72: res = 32'b00000000000000000011011110001101; // input=-0.265625, output=0.433981464804
            7'd73: res = 32'b00000000000000000011011010010010; // input=-0.296875, output=0.426321592547
            7'd74: res = 32'b00000000000000000011010110011000; // input=-0.328125, output=0.418696909356
            7'd75: res = 32'b00000000000000000011010010011111; // input=-0.359375, output=0.411110869232
            7'd76: res = 32'b00000000000000000011001110101000; // input=-0.390625, output=0.403566853735
            7'd77: res = 32'b00000000000000000011001010110010; // input=-0.421875, output=0.396068166274
            7'd78: res = 32'b00000000000000000011000110111110; // input=-0.453125, output=0.388618026706
            7'd79: res = 32'b00000000000000000011000011001100; // input=-0.484375, output=0.381219566256
            7'd80: res = 32'b00000000000000000010111111011011; // input=-0.515625, output=0.373875822772
            7'd81: res = 32'b00000000000000000010111011101100; // input=-0.546875, output=0.366589736322
            7'd82: res = 32'b00000000000000000010111000000000; // input=-0.578125, output=0.35936414516
            7'd83: res = 32'b00000000000000000010110100010101; // input=-0.609375, output=0.352201782048
            7'd84: res = 32'b00000000000000000010110000101100; // input=-0.640625, output=0.345105270958
            7'd85: res = 32'b00000000000000000010101101000110; // input=-0.671875, output=0.33807712415
            7'd86: res = 32'b00000000000000000010101001100010; // input=-0.703125, output=0.331119739629
            7'd87: res = 32'b00000000000000000010100110000001; // input=-0.734375, output=0.324235398981
            7'd88: res = 32'b00000000000000000010100010100001; // input=-0.765625, output=0.317426265588
            7'd89: res = 32'b00000000000000000010011111000101; // input=-0.796875, output=0.310694383215
            7'd90: res = 32'b00000000000000000010011011101011; // input=-0.828125, output=0.304041674967
            7'd91: res = 32'b00000000000000000010011000010011; // input=-0.859375, output=0.297469942605
            7'd92: res = 32'b00000000000000000010010100111111; // input=-0.890625, output=0.290980866215
            7'd93: res = 32'b00000000000000000010010001101101; // input=-0.921875, output=0.284576004217
            7'd94: res = 32'b00000000000000000010001110011110; // input=-0.953125, output=0.278256793702
            7'd95: res = 32'b00000000000000000010001011010010; // input=-0.984375, output=0.272024551094
            7'd96: res = 32'b00000000000000000010001000001000; // input=-1.015625, output=0.2658804731
            7'd97: res = 32'b00000000000000000010000101000010; // input=-1.046875, output=0.259825637961
            7'd98: res = 32'b00000000000000000010000001111111; // input=-1.078125, output=0.253861006969
            7'd99: res = 32'b00000000000000000001111110111110; // input=-1.109375, output=0.24798742624
            7'd100: res = 32'b00000000000000000001111100000001; // input=-1.140625, output=0.242205628725
            7'd101: res = 32'b00000000000000000001111001000110; // input=-1.171875, output=0.236516236446
            7'd102: res = 32'b00000000000000000001110110001111; // input=-1.203125, output=0.230919762929
            7'd103: res = 32'b00000000000000000001110011011010; // input=-1.234375, output=0.225416615835
            7'd104: res = 32'b00000000000000000001110000101001; // input=-1.265625, output=0.220007099746
            7'd105: res = 32'b00000000000000000001101101111011; // input=-1.296875, output=0.214691419112
            7'd106: res = 32'b00000000000000000001101011010000; // input=-1.328125, output=0.20946968133
            7'd107: res = 32'b00000000000000000001101000101000; // input=-1.359375, output=0.204341899937
            7'd108: res = 32'b00000000000000000001100110000011; // input=-1.390625, output=0.199307997904
            7'd109: res = 32'b00000000000000000001100011100001; // input=-1.421875, output=0.194367811019
            7'd110: res = 32'b00000000000000000001100001000010; // input=-1.453125, output=0.18952109133
            7'd111: res = 32'b00000000000000000001011110100110; // input=-1.484375, output=0.184767510648
            7'd112: res = 32'b00000000000000000001011100001110; // input=-1.515625, output=0.180106664086
            7'd113: res = 32'b00000000000000000001011001111000; // input=-1.546875, output=0.175538073623
            7'd114: res = 32'b00000000000000000001010111100101; // input=-1.578125, output=0.171061191679
            7'd115: res = 32'b00000000000000000001010101010110; // input=-1.609375, output=0.166675404688
            7'd116: res = 32'b00000000000000000001010011001001; // input=-1.640625, output=0.162380036667
            7'd117: res = 32'b00000000000000000001010000111111; // input=-1.671875, output=0.158174352748
            7'd118: res = 32'b00000000000000000001001110111000; // input=-1.703125, output=0.154057562691
            7'd119: res = 32'b00000000000000000001001100110100; // input=-1.734375, output=0.150028824342
            7'd120: res = 32'b00000000000000000001001010110011; // input=-1.765625, output=0.146087247048
            7'd121: res = 32'b00000000000000000001001000110101; // input=-1.796875, output=0.14223189501
            7'd122: res = 32'b00000000000000000001000110111001; // input=-1.828125, output=0.138461790569
            7'd123: res = 32'b00000000000000000001000101000000; // input=-1.859375, output=0.134775917423
            7'd124: res = 32'b00000000000000000001000011001010; // input=-1.890625, output=0.131173223762
            7'd125: res = 32'b00000000000000000001000001010111; // input=-1.921875, output=0.127652625322
            7'd126: res = 32'b00000000000000000000111111100110; // input=-1.953125, output=0.124213008352
            7'd127: res = 32'b00000000000000000000111101111000; // input=-1.984375, output=0.12085323249
        endcase
    end
    converter U0 (
        .a(in),
        .index(index)
    );

endmodule

module converter(a, index);
        input  [31:0] a;
        output [6:0] index;

        assign index[6] = a[31];
        assign index[5:5] = a[15:15];
        assign index[4:0] = a[14:10];
endmodule
