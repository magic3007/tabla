`timescale 1ns/1ps
module comp(
    in1,
    in2,
    out
);

	// *****************************************************************************
	parameter   LEN = 8;

	// *****************************************************************************
	input	[LEN - 1 : 0]   in1;
	input	[LEN - 1 : 0]   in2;
	output out;

	// *****************************************************************************
	assign out = ( in1 >= in2 ) ? 0 : 1;

endmodule
