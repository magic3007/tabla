module zynq_wrapper #(
    parameter READ_ADDR_BASE_0   = 32'h00000000,
    parameter WRITE_ADDR_BASE_0  = 32'h02000000
)
(
    inout wire [14:0]   DDR_addr,
    inout wire [2:0]    DDR_ba,
    inout wire          DDR_cas_n,
    inout wire          DDR_ck_n,
    inout wire          DDR_ck_p,
    inout wire          DDR_cke,
    inout wire          DDR_cs_n,
    inout wire [3:0]    DDR_dm,
    inout wire [31:0]   DDR_dq,
    inout wire [3:0]    DDR_dqs_n,
    inout wire [3:0]    DDR_dqs_p,
    inout wire          DDR_odt,
    inout wire          DDR_ras_n,
    inout wire          DDR_reset_n,
    inout wire          DDR_we_n,
    inout wire          FIXED_IO_ddr_vrn,
    inout wire          FIXED_IO_ddr_vrp,
    inout wire [53:0]   FIXED_IO_mio,
    inout wire          FIXED_IO_ps_clk,
    inout wire          FIXED_IO_ps_porb,
    inout wire          FIXED_IO_ps_srstb
    );

    wire                FCLK_CLK0;
    wire                FCLK_RESET0_N;

    wire [31:0]         M_AXI_GP0_awaddr;
    wire [2:0]          M_AXI_GP0_awprot;
    wire                M_AXI_GP0_awready;
    wire                M_AXI_GP0_awvalid;
    wire [31:0]         M_AXI_GP0_wdata;
    wire [3:0]          M_AXI_GP0_wstrb;
    wire                M_AXI_GP0_wvalid;
    wire                M_AXI_GP0_wready;
    wire [1:0]          M_AXI_GP0_bresp;
    wire                M_AXI_GP0_bvalid;
    wire                M_AXI_GP0_bready;
    wire [31:0]         M_AXI_GP0_araddr;
    wire [2:0]          M_AXI_GP0_arprot;
    wire                M_AXI_GP0_arvalid;
    wire                M_AXI_GP0_arready;
    wire [31:0]         M_AXI_GP0_rdata;
    wire [1:0]          M_AXI_GP0_rresp;
    wire                M_AXI_GP0_rvalid;
    wire                M_AXI_GP0_rready;

    wire [31:0]         S_AXI_HP0_araddr;
    wire [1:0]          S_AXI_HP0_arburst;
    wire [3:0]          S_AXI_HP0_arcache;
    wire [5:0]          S_AXI_HP0_arid;
    wire [3:0]          S_AXI_HP0_arlen;
    wire [1:0]          S_AXI_HP0_arlock;
    wire [2:0]          S_AXI_HP0_arprot;
    wire [3:0]          S_AXI_HP0_arqos;
    wire                S_AXI_HP0_arready;
    wire [2:0]          S_AXI_HP0_arsize;
    wire                S_AXI_HP0_arvalid;
    wire [31:0]         S_AXI_HP0_awaddr;
    wire [1:0]          S_AXI_HP0_awburst;
    wire [3:0]          S_AXI_HP0_awcache;
    wire [5:0]          S_AXI_HP0_awid;
    wire [3:0]          S_AXI_HP0_awlen;
    wire [1:0]          S_AXI_HP0_awlock;
    wire [2:0]          S_AXI_HP0_awprot;
    wire [3:0]          S_AXI_HP0_awqos;
    wire                S_AXI_HP0_awready;
    wire [2:0]          S_AXI_HP0_awsize;
    wire                S_AXI_HP0_awvalid;
    wire [5:0]          S_AXI_HP0_bid;
    wire                S_AXI_HP0_bready;
    wire [1:0]          S_AXI_HP0_bresp;
    wire                S_AXI_HP0_bvalid;
    wire [63:0]         S_AXI_HP0_rdata;
    wire [5:0]          S_AXI_HP0_rid;
    wire                S_AXI_HP0_rlast;
    wire                S_AXI_HP0_rready;
    wire [1:0]          S_AXI_HP0_rresp;
    wire                S_AXI_HP0_rvalid;
    wire [63:0]         S_AXI_HP0_wdata;
    wire [5:0]          S_AXI_HP0_wid;
    wire                S_AXI_HP0_wlast;
    wire                S_AXI_HP0_wready;
    wire [7:0]          S_AXI_HP0_wstrb;
    wire                S_AXI_HP0_wvalid;

    localparam integer  C_S_AXI_DATA_WIDTH    = 32;
    localparam integer  C_S_AXI_ADDR_WIDTH    = 32;
    localparam integer  C_M_AXI_DATA_WIDTH    = 64;
    localparam integer  C_M_AXI_ADDR_WIDTH    = 32;

    wire                                outBuf_empty;
    wire                                outBuf_pop;
    wire                                outBuf_full;
    wire                                outBuf_push;
    wire [FIFO_ADDR_WIDTH:0]            outBuf_count;
    wire [C_M_AXI_DATA_WIDTH-1:0]       data_to_outBuf;
    wire [C_M_AXI_DATA_WIDTH-1:0]       data_from_outBuf;
    wire                                inBuf_empty;
    wire                                inBuf_pop;
    wire                                inBuf_full;
    wire                                inBuf_push;
    wire [C_M_AXI_DATA_WIDTH-1:0]       data_to_inBuf;
    wire [C_M_AXI_DATA_WIDTH-1:0]       data_from_inBuf;
    wire [FIFO_ADDR_WIDTH:0]            inBuf_count;

    localparam integer FIFO_ADDR_WIDTH = 8;


    wire tx_req, tx_done;


  zynq zynq_i (
    .DDR_addr               ( DDR_addr            ),
    .DDR_ba                 ( DDR_ba              ),
    .DDR_cas_n              ( DDR_cas_n           ),
    .DDR_ck_n               ( DDR_ck_n            ),
    .DDR_ck_p               ( DDR_ck_p            ),
    .DDR_cke                ( DDR_cke             ),
    .DDR_cs_n               ( DDR_cs_n            ),
    .DDR_dm                 ( DDR_dm              ),
    .DDR_dq                 ( DDR_dq              ),
    .DDR_dqs_n              ( DDR_dqs_n           ),
    .DDR_dqs_p              ( DDR_dqs_p           ),
    .DDR_odt                ( DDR_odt             ),
    .DDR_ras_n              ( DDR_ras_n           ),
    .DDR_reset_n            ( DDR_reset_n         ),
    .DDR_we_n               ( DDR_we_n            ),

    .FIXED_IO_ddr_vrn       ( FIXED_IO_ddr_vrn    ),
    .FIXED_IO_ddr_vrp       ( FIXED_IO_ddr_vrp    ),
    .FIXED_IO_mio           ( FIXED_IO_mio        ),
    .FIXED_IO_ps_clk        ( FIXED_IO_ps_clk     ),
    .FIXED_IO_ps_porb       ( FIXED_IO_ps_porb    ),
    .FIXED_IO_ps_srstb      ( FIXED_IO_ps_srstb   ),

    .FCLK_CLK0              ( FCLK_CLK0           ),
    .FCLK_RESET0_N          ( FCLK_RESET0_N       ),

    .M_AXI_GP0_awaddr       ( M_AXI_GP0_awaddr    ),
    .M_AXI_GP0_awprot       ( M_AXI_GP0_awprot    ),
    .M_AXI_GP0_awready      ( M_AXI_GP0_awready   ),
    .M_AXI_GP0_awvalid      ( M_AXI_GP0_awvalid   ),
    .M_AXI_GP0_araddr       ( M_AXI_GP0_araddr    ),
    .M_AXI_GP0_arprot       ( M_AXI_GP0_arprot    ),
    .M_AXI_GP0_arready      ( M_AXI_GP0_arready   ),
    .M_AXI_GP0_arvalid      ( M_AXI_GP0_arvalid   ),
    .M_AXI_GP0_bready       ( M_AXI_GP0_bready    ),
    .M_AXI_GP0_bresp        ( M_AXI_GP0_bresp     ),
    .M_AXI_GP0_bvalid       ( M_AXI_GP0_bvalid    ),
    .M_AXI_GP0_rdata        ( M_AXI_GP0_rdata     ),
    .M_AXI_GP0_rready       ( M_AXI_GP0_rready    ),
    .M_AXI_GP0_rresp        ( M_AXI_GP0_rresp     ),
    .M_AXI_GP0_rvalid       ( M_AXI_GP0_rvalid    ),
    .M_AXI_GP0_wdata        ( M_AXI_GP0_wdata     ),
    .M_AXI_GP0_wready       ( M_AXI_GP0_wready    ),
    .M_AXI_GP0_wstrb        ( M_AXI_GP0_wstrb     ),
    .M_AXI_GP0_wvalid       ( M_AXI_GP0_wvalid    ),

    .S_AXI_HP0_araddr       ( S_AXI_HP0_araddr    ),
    .S_AXI_HP0_arburst      ( S_AXI_HP0_arburst   ),
    .S_AXI_HP0_arcache      ( S_AXI_HP0_arcache   ),
    .S_AXI_HP0_arid         ( S_AXI_HP0_arid      ),
    .S_AXI_HP0_arlen        ( S_AXI_HP0_arlen     ),
    .S_AXI_HP0_arlock       ( S_AXI_HP0_arlock    ),
    .S_AXI_HP0_arprot       ( S_AXI_HP0_arprot    ),
    .S_AXI_HP0_arqos        ( S_AXI_HP0_arqos     ),
    .S_AXI_HP0_arready      ( S_AXI_HP0_arready   ),
    .S_AXI_HP0_arsize       ( S_AXI_HP0_arsize    ),
    .S_AXI_HP0_arvalid      ( S_AXI_HP0_arvalid   ),
    .S_AXI_HP0_awaddr       ( S_AXI_HP0_awaddr    ),
    .S_AXI_HP0_awburst      ( S_AXI_HP0_awburst   ),
    .S_AXI_HP0_awcache      ( S_AXI_HP0_awcache   ),
    .S_AXI_HP0_awid         ( S_AXI_HP0_awid      ),
    .S_AXI_HP0_awlen        ( S_AXI_HP0_awlen     ),
    .S_AXI_HP0_awlock       ( S_AXI_HP0_awlock    ),
    .S_AXI_HP0_awprot       ( S_AXI_HP0_awprot    ),
    .S_AXI_HP0_awqos        ( S_AXI_HP0_awqos     ),
    .S_AXI_HP0_awready      ( S_AXI_HP0_awready   ),
    .S_AXI_HP0_awsize       ( S_AXI_HP0_awsize    ),
    .S_AXI_HP0_awvalid      ( S_AXI_HP0_awvalid   ),
    .S_AXI_HP0_bid          ( S_AXI_HP0_bid       ),
    .S_AXI_HP0_bready       ( S_AXI_HP0_bready    ),
    .S_AXI_HP0_bresp        ( S_AXI_HP0_bresp     ),
    .S_AXI_HP0_bvalid       ( S_AXI_HP0_bvalid    ),
    .S_AXI_HP0_rdata        ( S_AXI_HP0_rdata     ),
    .S_AXI_HP0_rid          ( S_AXI_HP0_rid       ),
    .S_AXI_HP0_rlast        ( S_AXI_HP0_rlast     ),
    .S_AXI_HP0_rready       ( S_AXI_HP0_rready    ),
    .S_AXI_HP0_rresp        ( S_AXI_HP0_rresp     ),
    .S_AXI_HP0_rvalid       ( S_AXI_HP0_rvalid    ),
    .S_AXI_HP0_wdata        ( S_AXI_HP0_wdata     ),
    //.S_AXI_HP0_wdata        ( 32'hAABACADA        ),
    .S_AXI_HP0_wid          ( S_AXI_HP0_wid       ),
    .S_AXI_HP0_wlast        ( S_AXI_HP0_wlast     ),
    .S_AXI_HP0_wready       ( S_AXI_HP0_wready    ),
    .S_AXI_HP0_wstrb        ( S_AXI_HP0_wstrb     ),
    .S_AXI_HP0_wvalid       ( S_AXI_HP0_wvalid    )
    );

axi_master #(
    .C_M_AXI_READ_TARGET    ( READ_ADDR_BASE_0    ),
    .C_M_AXI_WRITE_TARGET   ( WRITE_ADDR_BASE_0   )
) axim_hp0 (
    // System Signals
    .ACLK                   ( FCLK_CLK0           ),  //input
    .ARESETN                ( FCLK_RESET0_N       ),  //input
    
    // Master Interface Write Address
    .M_AXI_AWID             ( S_AXI_HP0_awid      ),  //output
    .M_AXI_AWADDR           ( S_AXI_HP0_awaddr    ),  //output
    .M_AXI_AWLEN            ( S_AXI_HP0_awlen     ),  //output
    .M_AXI_AWSIZE           ( S_AXI_HP0_awsize    ),  //output
    .M_AXI_AWBURST          ( S_AXI_HP0_awburst   ),  //output
    .M_AXI_AWLOCK           ( S_AXI_HP0_awlock    ),  //output
    .M_AXI_AWCACHE          ( S_AXI_HP0_awcache   ),  //output
    .M_AXI_AWPROT           ( S_AXI_HP0_awprot    ),  //output
    .M_AXI_AWQOS            ( S_AXI_HP0_awqos     ),  //output
    .M_AXI_AWVALID          ( S_AXI_HP0_awvalid   ),  //output
    .M_AXI_AWREADY          ( S_AXI_HP0_awready   ),  //input
    
    // Master Interface Write Data
    .M_AXI_WID              ( S_AXI_HP0_wid       ),  //output
    .M_AXI_WDATA            ( S_AXI_HP0_wdata     ),  //output
    .M_AXI_WSTRB            ( S_AXI_HP0_wstrb     ),  //output
    .M_AXI_WLAST            ( S_AXI_HP0_wlast     ),  //output
    .M_AXI_WVALID           ( S_AXI_HP0_wvalid    ),  //output
    .M_AXI_WREADY           ( S_AXI_HP0_wready    ),  //input
    
    // Master Interface Write Response
    .M_AXI_BID              ( S_AXI_HP0_bid       ),  //input
    .M_AXI_BRESP            ( S_AXI_HP0_bresp     ),  //input
    .M_AXI_BVALID           ( S_AXI_HP0_bvalid    ),  //input
    .M_AXI_BREADY           ( S_AXI_HP0_bready    ),  //output
   
    // Master Interface Read Address
    .M_AXI_ARID             ( S_AXI_HP0_arid      ),  //output
    .M_AXI_ARADDR           ( S_AXI_HP0_araddr    ),  //output
    .M_AXI_ARLEN            ( S_AXI_HP0_arlen     ),  //output
    .M_AXI_ARSIZE           ( S_AXI_HP0_arsize    ),  //output
    .M_AXI_ARBURST          ( S_AXI_HP0_arburst   ),  //output
    .M_AXI_ARLOCK           ( S_AXI_HP0_arlock    ),  //output
    .M_AXI_ARCACHE          ( S_AXI_HP0_arcache   ),  //output
    .M_AXI_ARQOS            ( S_AXI_HP0_arqos     ),  //output
    .M_AXI_ARPROT           ( S_AXI_HP0_arprot    ),  //output
    .M_AXI_ARVALID          ( S_AXI_HP0_arvalid   ),  //output
    .M_AXI_ARREADY          ( S_AXI_HP0_arready   ),  //input
    
    // Master Interface Read Data 
    .M_AXI_RID              ( S_AXI_HP0_rid       ),  //input
    .M_AXI_RDATA            ( S_AXI_HP0_rdata     ),  //input
    .M_AXI_RRESP            ( S_AXI_HP0_rresp     ),  //input
    .M_AXI_RLAST            ( S_AXI_HP0_rlast     ),  //input
    .M_AXI_RVALID           ( S_AXI_HP0_rvalid    ),  //input
    .M_AXI_RREADY           ( S_AXI_HP0_rready    ),  //output

    // NPU Design
    // WRITE from BRAM to DDR
    .outBuf_empty           ( outBuf_empty        ), //input
    .outBuf_pop             ( outBuf_pop          ), //output
    .data_from_outBuf       ( data_from_outBuf    ), //input
    //.data_from_outBuf       ( {16'hAAAA, data_from_outBuf[47:32], 16'hAAAA, data_from_outBuf[15:0]} ), //input
    .outBuf_count           ( outBuf_count        ), //input

    // READ from DDR to BRAM
    .data_to_inBuf          ( data_to_inBuf       ), //output
    .inBuf_push             ( inBuf_push          ), //output
    .inBuf_full             ( inBuf_full          ), //input
    .inBuf_count            ( inBuf_count         ), //input

    .tx_req                 ( tx_req              ), //input
    .tx_done                ( tx_done             )  //output
    ); 

fifo #(
    .DATA_WIDTH             ( 64                  ),
    .ADDR_WIDTH             ( FIFO_ADDR_WIDTH     )
) fifo_inBuf (
    .clk                    ( FCLK_CLK0           ), //input
    .reset                  ( !FCLK_RESET0_N      ), //input
    .push                   ( inBuf_push          ), //input
    .pop                    ( inBuf_pop           ), //input
    .data_in                ( data_to_inBuf       ), //input
    .data_out               ( data_from_inBuf     ), //output
    .empty                  ( inBuf_empty         ), //output
    .full                   ( inBuf_full          ), //output
    .fifo_count             ( inBuf_count         )  //output
);

accelerator #(
    .DATA_WIDTH             ( 64                  ),
    .BUFFER_ADDR_WIDTH      ( FIFO_ADDR_WIDTH     ),
    .TYPE                   ( "LOOPBACK"        )
) tabla (
    .ACLK                   ( FCLK_CLK0           ), //input
    .ARESETN                ( FCLK_RESET0_N       ), //input
    .inBuf_empty            ( inBuf_empty         ), //input
    .inBuf_count            ( inBuf_count         ), //input
    .inBuf_pop              ( inBuf_pop           ), //output
    .data_from_inBuf        ( data_from_inBuf     ), //input
    .outBuf_full            ( outBuf_full         ), //input
    .outBuf_count           ( outBuf_count        ), //input
    .outBuf_push            ( outBuf_push         ), //output
    .data_to_outBuf         ( data_to_outBuf      )  //output
);

fifo_fwft #(
    .DATA_WIDTH             ( 64                  ),
    .ADDR_WIDTH             ( FIFO_ADDR_WIDTH     )
) fifo_outBuf (
    .clk                    ( FCLK_CLK0           ),  //input
    .reset                  ( !FCLK_RESET0_N      ),  //input
    .push                   ( outBuf_push         ),  //input
    .pop                    ( outBuf_pop          ),  //input
    .data_in                ( data_to_outBuf      ),  //input
    .data_out               ( data_from_outBuf    ),  //output
    .empty                  ( outBuf_empty        ),  //output
    .full                   ( outBuf_full         ),  //output
    .fifo_count             ( outBuf_count        )   //output
);

axi4lite_slave #(
    .C_S_AXI_DATA_WIDTH     ( C_S_AXI_DATA_WIDTH  ),
    .C_S_AXI_ADDR_WIDTH     ( C_S_AXI_ADDR_WIDTH  )
) axi_slave_i (
    .S_AXI_ACLK             ( FCLK_CLK0           ),  //input
    .S_AXI_ARESETN          ( FCLK_RESET0_N       ),  //input

    .S_AXI_AWADDR           ( M_AXI_GP0_awaddr    ),  //input
    .S_AXI_AWPROT           ( M_AXI_GP0_awprot    ),  //input
    .S_AXI_AWVALID          ( M_AXI_GP0_awvalid   ),  //input
    .S_AXI_AWREADY          ( M_AXI_GP0_awready   ),  //output

    .S_AXI_WDATA            ( M_AXI_GP0_wdata     ),  //input
    .S_AXI_WSTRB            ( M_AXI_GP0_wstrb     ),  //input
    .S_AXI_WVALID           ( M_AXI_GP0_wvalid    ),  //input
    .S_AXI_WREADY           ( M_AXI_GP0_wready    ),  //output

    .S_AXI_BRESP            ( M_AXI_GP0_bresp     ),  //output
    .S_AXI_BVALID           ( M_AXI_GP0_bvalid    ),  //output
    .S_AXI_BREADY           ( M_AXI_GP0_bready    ),  //input

    .S_AXI_ARADDR           ( M_AXI_GP0_araddr    ),  //input
    .S_AXI_ARPROT           ( M_AXI_GP0_arprot    ),  //input
    .S_AXI_ARVALID          ( M_AXI_GP0_arvalid   ),  //input
    .S_AXI_ARREADY          ( M_AXI_GP0_arready   ),  //output

    .S_AXI_RDATA            ( M_AXI_GP0_rdata     ),  //output
    .S_AXI_RRESP            ( M_AXI_GP0_rresp     ),  //output
    .S_AXI_RVALID           ( M_AXI_GP0_rvalid    ),  //output
    .S_AXI_RREADY           ( M_AXI_GP0_rready    ),  //input

    .tx_req                 ( tx_req              ),  //output
    .tx_done                ( tx_done             )   //input
);

endmodule
